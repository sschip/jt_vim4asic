// module definition
module_000 u_module(
);

module_001 u_module();

module_002 
u_module();

module_003 
u_module
();

module_004 #(.PARAM_000(100))
u_module
();
// class definition
class_000 class_inst;
// task definition
// function definition
