// module definition
module module_000(
);

module module_001();

module 
module_002();

module 
module_003
();

module #(parameter PARAM_000 = 100)
module_004
();
// class definition
class class_000;
endclass
// task definition
// function definition
function uvm_component uvm_compnent::function_000 (string requested_type_name,
                                                       string name);
                                                   return factory.create_component_by_name(requested_type_name, get_full_name(),
                                                                                           name, this);
endfunction
